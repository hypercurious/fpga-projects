module bin_2_7 (x, s);
    input  [3:0] x;
    output [6:0] s;
  
    assign s = (x == 4'd0 ) ? 7'b1111110 :
               (x == 4'd1 ) ? 7'b0110000 :
               (x == 4'd2 ) ? 7'b1101101 :
               (x == 4'd3 ) ? 7'b1111001 :
               (x == 4'd4 ) ? 7'b0110011 :
               (x == 4'd5 ) ? 7'b1011011 :
               (x == 4'd6 ) ? 7'b1011111 :
               (x == 4'd7 ) ? 7'b1110010 :
               (x == 4'd8 ) ? 7'b1111111 :
               (x == 4'd9 ) ? 7'b1111011 :
               (x == 4'd10) ? 7'b1110111 :
               (x == 4'd11) ? 7'b0011111 :
               (x == 4'd12) ? 7'b1001110 :
               (x == 4'd13) ? 7'b0111101 :
               (x == 4'd14) ? 7'b1001111 : 7'b1000111 ;
endmodule
             
