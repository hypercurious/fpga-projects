module ask6_2a(a,b,s);
    input [1:0]a,b;
    output reg [6:0]s;
    wire [3:0]o;
    
    assign o = a*b;
    
    always @ (o) begin
        case(o)
            4'b0000:
                 s[6:0]=7'b1110111;
            4'b0001:
                 s[6:0]=7'b0010010;
            4'b0010:
                 s[6:0]=7'b1011101;
            4'b0011:
                 s[6:0]=7'b1011011;
            4'b0100:
                 s[6:0]=7'b0111010;
            4'b0101:
                 s[6:0]=7'b1101011;
            4'b0110:
                 s[6:0]=7'b1101111;
            4'b0111:
                 s[6:0]=7'b1010010;
            4'b1000:
                 s[6:0]=7'b1111111;
            4'b1001:
                 s[6:0]=7'b1111011;
            default:
                 s[6:0]=7'b0000000;
        endcase
    end
    
endmodule
