library verilog;
use verilog.vl_types.all;
entity testcounter_8bit is
end testcounter_8bit;
