module bin_2_led (x,s);
    input  [3:0] x;
    output [9:0] s;
    
    assign s = (x == 4'd0 ) ? 10'b0000000000 :
               (x == 4'd1 ) ? 10'b0000000001 :
               (x == 4'd2 ) ? 10'b0000000011 :
               (x == 4'd3 ) ? 10'b0000000111 :
               (x == 4'd4 ) ? 10'b0000001111 :
               (x == 4'd5 ) ? 10'b0000011111 :
               (x == 4'd6 ) ? 10'b0000111111 :
               (x == 4'd7 ) ? 10'b0001111111 :
               (x == 4'd8 ) ? 10'b0011111111 :
               (x == 4'd9 ) ? 10'b0111111111 :
               (x == 4'd10) ? 10'b1111111111 : 10'b0101010101 ;
endmodule
