library verilog;
use verilog.vl_types.all;
entity test_sync_counter_8bit is
end test_sync_counter_8bit;
